// Module: when buttons 1 and 2 are pressed, turn on LED
module and_gate (
